        rom[255] = 8'b01001000;
        rom[254] = 8'b11000001;
        rom[253] = 8'b00111000;
        rom[252] = 8'b00111110;
        rom[251] = 8'b10111100;
        rom[250] = 8'b01001100;
        rom[249] = 8'b01100101;
        rom[248] = 8'b00010011;
        rom[247] = 8'b01101010;
        rom[246] = 8'b11011011;
        rom[245] = 8'b00010010;
        rom[244] = 8'b11011111;
        rom[243] = 8'b11101111;
        rom[242] = 8'b11100111;
        rom[241] = 8'b10001111;
        rom[240] = 8'b00110111;
        rom[239] = 8'b11001100;
        rom[238] = 8'b01010110;
        rom[237] = 8'b10111001;
        rom[236] = 8'b00100011;
        rom[235] = 8'b11011110;
        rom[234] = 8'b10010010;
        rom[233] = 8'b10101001;
        rom[232] = 8'b11100111;
        rom[231] = 8'b00001101;
        rom[230] = 8'b10111110;
        rom[229] = 8'b10100010;
        rom[228] = 8'b11100011;
        rom[227] = 8'b01100100;
        rom[226] = 8'b01101010;
        rom[225] = 8'b00100011;
        rom[224] = 8'b11011010;
        rom[223] = 8'b01111110;
        rom[222] = 8'b00110000;
        rom[221] = 8'b01100011;
        rom[220] = 8'b11100001;
        rom[219] = 8'b10000010;
        rom[218] = 8'b10010001;
        rom[217] = 8'b00111011;
        rom[216] = 8'b01100000;
        rom[215] = 8'b11110001;
        rom[214] = 8'b01110000;
        rom[213] = 8'b01001111;
        rom[212] = 8'b00001110;
        rom[211] = 8'b00100110;
        rom[210] = 8'b11111000;
        rom[209] = 8'b00001011;
        rom[208] = 8'b00010000;
        rom[207] = 8'b01001010;
        rom[206] = 8'b10011110;
        rom[205] = 8'b11100011;
        rom[204] = 8'b10011011;
        rom[203] = 8'b11110110;
        rom[202] = 8'b00110011;
        rom[201] = 8'b11010110;
        rom[200] = 8'b01001110;
        rom[199] = 8'b10101000;
        rom[198] = 8'b01100001;
        rom[197] = 8'b11100000;
        rom[196] = 8'b00101111;
        rom[195] = 8'b11110100;
        rom[194] = 8'b00111000;
        rom[193] = 8'b11011101;
        rom[192] = 8'b11111010;
        rom[191] = 8'b00000100;
        rom[190] = 8'b01101001;
        rom[189] = 8'b00111101;
        rom[188] = 8'b10101110;
        rom[187] = 8'b11111100;
        rom[186] = 8'b10100111;
        rom[185] = 8'b11100101;
        rom[184] = 8'b10001100;
        rom[183] = 8'b11100010;
        rom[182] = 8'b00110101;
        rom[181] = 8'b11100111;
        rom[180] = 8'b11010111;
        rom[179] = 8'b11101010;
        rom[178] = 8'b00000111;
        rom[177] = 8'b10011100;
        rom[176] = 8'b01110111;
        rom[175] = 8'b11100100;
        rom[174] = 8'b01110000;
        rom[173] = 8'b00111100;
        rom[172] = 8'b11011100;
        rom[171] = 8'b00100101;
        rom[170] = 8'b01100000;
        rom[169] = 8'b10110000;
        rom[168] = 8'b01010000;
        rom[167] = 8'b01101110;
        rom[166] = 8'b10011101;
        rom[165] = 8'b00010111;
        rom[164] = 8'b01001100;
        rom[163] = 8'b11010001;
        rom[162] = 8'b10101001;
        rom[161] = 8'b00111111;
        rom[160] = 8'b11111100;
        rom[159] = 8'b11100011;
        rom[158] = 8'b10000111;
        rom[157] = 8'b11101101;
        rom[156] = 8'b10001011;
        rom[155] = 8'b01000100;
        rom[154] = 8'b00111000;
        rom[153] = 8'b11110010;
        rom[152] = 8'b00011111;
        rom[151] = 8'b10000010;
        rom[150] = 8'b00011000;
        rom[149] = 8'b10100100;
        rom[148] = 8'b01100000;
        rom[147] = 8'b01101101;
        rom[146] = 8'b11100100;
        rom[145] = 8'b10101001;
        rom[144] = 8'b01001000;
        rom[143] = 8'b01001001;
        rom[142] = 8'b10010011;
        rom[141] = 8'b10110011;
        rom[140] = 8'b01110100;
        rom[139] = 8'b10011000;
        rom[138] = 8'b00101000;
        rom[137] = 8'b11101001;
        rom[136] = 8'b10001000;
        rom[135] = 8'b01011100;
        rom[134] = 8'b01010000;
        rom[133] = 8'b01101111;
        rom[132] = 8'b11010010;
        rom[131] = 8'b01111001;
        rom[130] = 8'b11100110;
        rom[129] = 8'b10000110;
        rom[128] = 8'b11101011;
        rom[127] = 8'b10001001;
        rom[126] = 8'b00110011;
        rom[125] = 8'b01010111;
        rom[124] = 8'b11101010;
        rom[123] = 8'b10110101;
        rom[122] = 8'b01010010;
        rom[121] = 8'b10110100;
        rom[120] = 8'b00001001;
        rom[119] = 8'b00110000;
        rom[118] = 8'b10000100;
        rom[117] = 8'b00010001;
        rom[116] = 8'b10011001;
        rom[115] = 8'b11000100;
        rom[114] = 8'b11100001;
        rom[113] = 8'b01001010;
        rom[112] = 8'b00110101;
        rom[111] = 8'b10000001;
        rom[110] = 8'b10111100;
        rom[109] = 8'b11100100;
        rom[108] = 8'b01010100;
        rom[107] = 8'b00101111;
        rom[106] = 8'b10000101;
        rom[105] = 8'b10011001;
        rom[104] = 8'b00100101;
        rom[103] = 8'b10110001;
        rom[102] = 8'b01010101;
        rom[101] = 8'b00000001;
        rom[100] = 8'b11100110;
        rom[ 99] = 8'b11001000;
        rom[ 98] = 8'b10111011;
        rom[ 97] = 8'b00111000;
        rom[ 96] = 8'b00000001;
        rom[ 95] = 8'b11101011;
        rom[ 94] = 8'b00111011;
        rom[ 93] = 8'b11011100;
        rom[ 92] = 8'b11001100;
        rom[ 91] = 8'b11100000;
        rom[ 90] = 8'b01111010;
        rom[ 89] = 8'b10001001;
        rom[ 88] = 8'b00011110;
        rom[ 87] = 8'b00110001;
        rom[ 86] = 8'b01001110;
        rom[ 85] = 8'b10110001;
        rom[ 84] = 8'b01011010;
        rom[ 83] = 8'b00100001;
        rom[ 82] = 8'b11110111;
        rom[ 81] = 8'b11101101;
        rom[ 80] = 8'b11000001;
        rom[ 79] = 8'b11101011;
        rom[ 78] = 8'b01000111;
        rom[ 77] = 8'b10101001;
        rom[ 76] = 8'b11011111;
        rom[ 75] = 8'b00000110;
        rom[ 74] = 8'b10111011;
        rom[ 73] = 8'b01101101;
        rom[ 72] = 8'b00110011;
        rom[ 71] = 8'b11101011;
        rom[ 70] = 8'b10010101;
        rom[ 69] = 8'b01001100;
        rom[ 68] = 8'b11110001;
        rom[ 67] = 8'b11000111;
        rom[ 66] = 8'b01000111;
        rom[ 65] = 8'b00011110;
        rom[ 64] = 8'b11011100;
        rom[ 63] = 8'b11010101;
        rom[ 62] = 8'b11011111;
        rom[ 61] = 8'b01100011;
        rom[ 60] = 8'b00001001;
        rom[ 59] = 8'b11010110;
        rom[ 58] = 8'b00111111;
        rom[ 57] = 8'b10101010;
        rom[ 56] = 8'b11101111;
        rom[ 55] = 8'b11011000;
        rom[ 54] = 8'b01000000;
        rom[ 53] = 8'b00111010;
        rom[ 52] = 8'b00000111;
        rom[ 51] = 8'b11101001;
        rom[ 50] = 8'b10111001;
        rom[ 49] = 8'b01000011;
        rom[ 48] = 8'b00101001;
        rom[ 47] = 8'b10001010;
        rom[ 46] = 8'b01111110;
        rom[ 45] = 8'b01110010;
        rom[ 44] = 8'b00110010;
        rom[ 43] = 8'b11111011;
        rom[ 42] = 8'b00111111;
        rom[ 41] = 8'b11010000;
        rom[ 40] = 8'b00111111;
        rom[ 39] = 8'b01011001;
        rom[ 38] = 8'b01011001;
        rom[ 37] = 8'b10101101;
        rom[ 36] = 8'b00010101;
        rom[ 35] = 8'b01010000;
        rom[ 34] = 8'b01111101;
        rom[ 33] = 8'b01001111;
        rom[ 32] = 8'b00111100;
        rom[ 31] = 8'b10000000;
        rom[ 30] = 8'b00100011;
        rom[ 29] = 8'b01011101;
        rom[ 28] = 8'b00000100;
        rom[ 27] = 8'b10001001;
        rom[ 26] = 8'b10001001;
        rom[ 25] = 8'b01101001;
        rom[ 24] = 8'b01011011;
        rom[ 23] = 8'b10101001;
        rom[ 22] = 8'b01111111;
        rom[ 21] = 8'b11100111;
        rom[ 20] = 8'b10010110;
        rom[ 19] = 8'b10111111;
        rom[ 18] = 8'b00111010;
        rom[ 17] = 8'b00010010;
        rom[ 16] = 8'b00000010;
        rom[ 15] = 8'b11011001;
        rom[ 14] = 8'b01101111;
        rom[ 13] = 8'b11110000;
        rom[ 12] = 8'b11101100;
        rom[ 11] = 8'b10010010;
        rom[ 10] = 8'b10110011;
        rom[  9] = 8'b01001011;
        rom[  8] = 8'b11010100;
        rom[  7] = 8'b00001110;
        rom[  6] = 8'b01000000;
        rom[  5] = 8'b01111111;
        rom[  4] = 8'b11000011;
        rom[  3] = 8'b10100110;
        rom[  2] = 8'b01111000;
        rom[  1] = 8'b01000100;
        rom[  0] = 8'b01001011;
