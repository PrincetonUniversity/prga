module fifo_tb();
endmodule