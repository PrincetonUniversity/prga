//# 3 inputs
//# 6 outputs
//# 21 D-type flipflops
//# 59 inverters
//# 99 gates (11 ANDs + 30 NANDs + 24 ORs + 34 NORs)

module s382(clk,CLR,FM,GRN1,GRN2,RED1,RED2,TEST,YLW1,YLW2);
input clk,FM,TEST,CLR;
output GRN1,GRN2,RED1,YLW2,RED2,YLW1;

  wire TESTL,TESTLVIINLATCHVCDAD,FML,FMLVIINLATCHVCDAD,OLATCH_Y2L,TCOMB_YA2,
    OLATCHVUC_6,Y1C,OLATCHVUC_5,R2C,OLATCH_R1L,TCOMB_RA1,OLATCH_G2L,TCOMB_GA2,
    OLATCH_G1L,TCOMB_GA1,OLATCH_FEL,TCOMB_FE_BF,C3_Q3,C3_Q3VD,C3_Q2,C3_Q2VD,
    C3_Q1,C3_Q1VD,C3_Q0,C3_Q0VD,UC_16,UC_16VD,UC_17,UC_17VD,UC_18,UC_18VD,
    UC_19,UC_19VD,UC_8,UC_8VD,UC_9,UC_9VD,UC_10,UC_10VD,UC_11,UC_11VD,
    TESTLVIINLATCHN,FMLVIINLATCHN,OLATCH_Y1L,OLATCH_R2L,UC_23,UC_24,UC_25,
    UC_26,UC_20,C2_QN2,UC_21,UC_22,UC_12,UC_13,UC_14,UC_15,FMBVIIR1,CLRBVIIR1,
    TCOMBVNFM,TESTBVIIR1,TCOMBVNQA,TCOMBVNQB,TCOMBVNQC,TCOMBVNQD,UC_11VUC_0,
    OUTBUFVBUFG1VIIR1,OUTBUFVBUFG2VIIR1,TCOMBVNFEL,OUTBUFVBUFR1VIIR1,
    OUTBUFVBUFY2VIIR1,FMB,CLRB,TESTB,UC_11VZ,C1VCO0,OUTBUFVBUFR2VIIR1,
    OUTBUFVBUFY1VIIR1,FMLVIINMUXVIIR1,TESTLVIINLATCHVCDN,FMLVIINLATCHVCDN,
    TCOMBVNCLR,TESTLVIINMUXVIIR1,C2VIINHN,CTST,UC_8VZ,UC_8VZVOR1NF,CO2,C2_CO,
    FMLVIINMUX,FMLVIINMUXVND1,TESTLVIINMUX,TESTLVIINMUXVND1,II84,TCOMB_FE,FEN,
    UC_16VZ,UC_16VZVOR1NF,C3VIINHN,C3_Q3VZ,C3_Q3VZVOR1NF,TCOMB_GA1VAD1NF,
    TCOMBVNODE6,TCOMB_GA2VAD4NF,TCOMB_GA2VAD3NF,TCOMB_GA2VAD2NF,
    TCOMB_GA2VAD1NF,R2CVAD1NF,Y1CVAD1NF,TCOMB_YA1,Y1CVAD2NF,R2CVAD2NF,
    TCOMB_RA2,TCOMB_RA1VOR2NF,TCOMBVNODE8VOR1NF,TCOMB_RA1VOR1NF,
    TCOMBVNODE8VOR2NF,FMLVIINMUXVOR1NF,TCOMB_RA2VOR3NF,TCOMB_RA2VOR1NF,
    TCOMBVNODE4VOR2NF,TCOMBVNODE4VOR1NF,TESTLVIINMUXVOR1NF,TCOMBVNODE16VOR1NF,
    TCOMBVNODE18,C1VCO2,UC_9VZVOR1NF,C1VCO1,UC_10VZVOR1NF,FMLVIINMUXVOR2NF,
    TESTLVIINMUXVOR2NF,C2VCO2,UC_17VZVOR1NF,C2VCO1,UC_18VZVOR1NF,C2VCO0,
    UC_19VZVOR1NF,C3VCO2,C3_Q2VZVOR1NF,C3VCO1,C3_Q1VZVOR1NF,C3VCO0,
    C3_Q0VZVOR1NF,UC_9VUC_0,UC_10VUC_0,TCOMBVNODE4,TCOMBVNODE14,TCOMBVNODE15,
    TCOMBVNODE12,TCOMBVNODE8,TCOMBVNODE16,TCOMBVNODE19,UC_9VZ,UC_10VZ,
    TCOMBVNODE3,UC_17VUC_0,UC_18VUC_0,UC_19VUC_0,UC_17VZ,UC_18VZ,UC_19VZ,
    C3_Q2VUC_0,C3_Q1VUC_0,C3_Q0VUC_0,C3_Q2VZ,C3_Q1VZ,C3_Q0VZ,C3VCIIA,C1VCIIA,
    C2VCIIA,C1_CO,UC_27;

  dff DFF_0(clk,TESTL,TESTLVIINLATCHVCDAD);
  dff DFF_1(clk,FML,FMLVIINLATCHVCDAD);
  dff DFF_2(clk,OLATCH_Y2L,TCOMB_YA2);
  dff DFF_3(clk,OLATCHVUC_6,Y1C);
  dff DFF_4(clk,OLATCHVUC_5,R2C);
  dff DFF_5(clk,OLATCH_R1L,TCOMB_RA1);
  dff DFF_6(clk,OLATCH_G2L,TCOMB_GA2);
  dff DFF_7(clk,OLATCH_G1L,TCOMB_GA1);
  dff DFF_8(clk,OLATCH_FEL,TCOMB_FE_BF);
  dff DFF_9(clk,C3_Q3,C3_Q3VD);
  dff DFF_10(clk,C3_Q2,C3_Q2VD);
  dff DFF_11(clk,C3_Q1,C3_Q1VD);
  dff DFF_12(clk,C3_Q0,C3_Q0VD);
  dff DFF_13(clk,UC_16,UC_16VD);
  dff DFF_14(clk,UC_17,UC_17VD);
  dff DFF_15(clk,UC_18,UC_18VD);
  dff DFF_16(clk,UC_19,UC_19VD);
  dff DFF_17(clk,UC_8,UC_8VD);
  dff DFF_18(clk,UC_9,UC_9VD);
  dff DFF_19(clk,UC_10,UC_10VD);
  dff DFF_20(clk,UC_11,UC_11VD);
  not NOT_0(TESTLVIINLATCHN,TESTL);
  not NOT_1(FMLVIINLATCHN,FML);
  not NOT_2(OLATCH_Y1L,OLATCHVUC_6);
  not NOT_3(OLATCH_R2L,OLATCHVUC_5);
  not NOT_4(UC_23,C3_Q3);
  not NOT_5(UC_24,C3_Q2);
  not NOT_6(UC_25,C3_Q1);
  not NOT_7(UC_26,C3_Q0);
  not NOT_8(UC_20,UC_16);
  not NOT_9(C2_QN2,UC_17);
  not NOT_10(UC_21,UC_18);
  not NOT_11(UC_22,UC_19);
  not NOT_12(UC_12,UC_8);
  not NOT_13(UC_13,UC_9);
  not NOT_14(UC_14,UC_10);
  not NOT_15(UC_15,UC_11);
  not NOT_16(FMBVIIR1,FM);
  not NOT_17(CLRBVIIR1,CLR);
  not NOT_18(TCOMBVNFM,FML);
  not NOT_19(TESTBVIIR1,TEST);
  not NOT_20(TCOMBVNQA,C3_Q0);
  not NOT_21(TCOMBVNQB,C3_Q1);
  not NOT_22(TCOMBVNQC,C3_Q2);
  not NOT_23(TCOMBVNQD,C3_Q3);
  not NOT_24(UC_11VUC_0,UC_11);
  not NOT_25(OUTBUFVBUFG1VIIR1,OLATCH_G1L);
  not NOT_26(OUTBUFVBUFG2VIIR1,OLATCH_G2L);
  not NOT_27(TCOMBVNFEL,OLATCH_FEL);
  not NOT_28(OUTBUFVBUFR1VIIR1,OLATCH_R1L);
  not NOT_29(OUTBUFVBUFY2VIIR1,OLATCH_Y2L);
  not NOT_30(FMB,FMBVIIR1);
  not NOT_31(CLRB,CLRBVIIR1);
  not NOT_32(TESTB,TESTBVIIR1);
  not NOT_33(UC_11VZ,UC_11VUC_0);
  not NOT_34(C1VCO0,UC_15);
  not NOT_35(GRN1,OUTBUFVBUFG1VIIR1);
  not NOT_36(GRN2,OUTBUFVBUFG2VIIR1);
  not NOT_37(RED1,OUTBUFVBUFR1VIIR1);
  not NOT_38(YLW2,OUTBUFVBUFY2VIIR1);
  not NOT_39(OUTBUFVBUFR2VIIR1,OLATCH_R2L);
  not NOT_40(OUTBUFVBUFY1VIIR1,OLATCH_Y1L);
  not NOT_41(FMLVIINMUXVIIR1,FMB);
  not NOT_42(TESTLVIINLATCHVCDN,CLRB);
  not NOT_43(FMLVIINLATCHVCDN,CLRB);
  not NOT_44(TCOMBVNCLR,CLRB);
  not NOT_45(TESTLVIINMUXVIIR1,TESTB);
  not NOT_46(RED2,OUTBUFVBUFR2VIIR1);
  not NOT_47(YLW1,OUTBUFVBUFY1VIIR1);
  not NOT_48(C2VIINHN,CTST);
  not NOT_49(UC_8VZ,UC_8VZVOR1NF);
  not NOT_50(CO2,C2_CO);
  not NOT_51(FMLVIINMUX,FMLVIINMUXVND1);
  not NOT_52(TESTLVIINMUX,TESTLVIINMUXVND1);
  not NOT_53(II84,TCOMB_FE);
  not NOT_54(FEN,TCOMB_FE);
  not NOT_55(UC_16VZ,UC_16VZVOR1NF);
  not NOT_56(C3VIINHN,CO2);
  not NOT_57(TCOMB_FE_BF,II84);
  not NOT_58(C3_Q3VZ,C3_Q3VZVOR1NF);
  and AND2_0(TCOMB_GA1VAD1NF,TCOMBVNODE6,OLATCH_FEL);
  and AND2_1(TCOMB_GA2VAD4NF,OLATCH_FEL,TCOMBVNCLR);
  and AND2_2(TCOMB_GA2VAD3NF,C3_Q2,TCOMBVNCLR);
  and AND3_0(TCOMB_GA2VAD2NF,C3_Q0,C3_Q1,TCOMBVNCLR);
  and AND3_1(TCOMB_GA2VAD1NF,TCOMBVNQA,C3_Q3,TCOMBVNCLR);
  and AND2_3(R2CVAD1NF,TCOMB_FE,C2_QN2);
  and AND2_4(FMLVIINLATCHVCDAD,FMLVIINLATCHVCDN,FMLVIINMUX);
  and AND2_5(Y1CVAD1NF,TCOMB_YA1,C2_QN2);
  and AND2_6(TESTLVIINLATCHVCDAD,TESTLVIINLATCHVCDN,TESTLVIINMUX);
  and AND2_7(Y1CVAD2NF,FEN,TCOMB_YA1);
  and AND2_8(R2CVAD2NF,FEN,TCOMB_RA2);
  or OR3_0(TCOMB_RA1VOR2NF,C3_Q2,C3_Q3,OLATCH_FEL);
  or OR3_1(TCOMBVNODE8VOR1NF,C3_Q0,C3_Q1,TCOMBVNFM);
  or OR4_0(TCOMB_RA1VOR1NF,TCOMBVNQA,C3_Q1,C3_Q2,OLATCH_FEL);
  or OR2_0(TCOMBVNODE8VOR2NF,TCOMBVNQD,TCOMBVNFM);
  or OR2_1(FMLVIINMUXVOR1NF,FMB,FML);
  or OR2_2(TCOMB_RA2VOR3NF,TCOMBVNQC,CLRB);
  or OR4_1(TCOMB_RA2VOR1NF,C3_Q0,C3_Q1,TCOMBVNQD,CLRB);
  or OR3_2(TCOMBVNODE4VOR2NF,C3_Q2,TCOMBVNQD,CLRB);
  or OR4_2(TCOMBVNODE4VOR1NF,TCOMBVNQC,C3_Q3,TCOMBVNFM,CLRB);
  or OR2_3(TESTLVIINMUXVOR1NF,TESTB,TESTL);
  or OR4_3(TCOMBVNODE16VOR1NF,TCOMBVNODE18,FML,C3_Q3,TCOMBVNQC);
  or OR2_4(UC_8VZVOR1NF,C1VCO2,UC_8);
  or OR2_5(UC_9VZVOR1NF,C1VCO1,UC_9);
  or OR2_6(UC_10VZVOR1NF,C1VCO0,UC_10);
  or OR2_7(FMLVIINMUXVOR2NF,FMLVIINMUXVIIR1,FMLVIINLATCHN);
  or OR2_8(TESTLVIINMUXVOR2NF,TESTLVIINMUXVIIR1,TESTLVIINLATCHN);
  or OR2_9(UC_16VZVOR1NF,C2VCO2,UC_16);
  or OR2_10(UC_17VZVOR1NF,C2VCO1,UC_17);
  or OR2_11(UC_18VZVOR1NF,C2VCO0,UC_18);
  or OR2_12(UC_19VZVOR1NF,C2VIINHN,UC_19);
  or OR2_13(C3_Q3VZVOR1NF,C3VCO2,C3_Q3);
  or OR2_14(C3_Q2VZVOR1NF,C3VCO1,C3_Q2);
  or OR2_15(C3_Q1VZVOR1NF,C3VCO0,C3_Q1);
  or OR2_16(C3_Q0VZVOR1NF,C3VIINHN,C3_Q0);
  nand NAND2_0(TCOMBVNODE18,TCOMBVNQB,C3_Q0);
  nand NAND4_0(TCOMBVNODE6,TCOMBVNFM,TCOMBVNQD,TCOMBVNQB,C3_Q0);
  nand NAND2_1(UC_9VUC_0,C1VCO1,UC_9);
  nand NAND2_2(UC_10VUC_0,C1VCO0,UC_10);
  nand NAND2_3(TCOMB_RA2,TCOMB_RA2VOR3NF,TCOMB_RA2VOR1NF);
  nand NAND2_4(TCOMBVNODE4,TCOMBVNODE4VOR2NF,TCOMBVNODE4VOR1NF);
  nand NAND2_5(TCOMBVNODE14,TCOMBVNODE15,TCOMBVNQA);
  nand NAND4_1(TCOMBVNODE12,TCOMBVNCLR,TCOMBVNFEL,TCOMBVNQC,C3_Q1);
  nand NAND4_2(TCOMBVNODE8,TCOMBVNCLR,C3_Q2,TCOMBVNODE8VOR2NF,
    TCOMBVNODE8VOR1NF);
  nand NAND3_0(TCOMB_RA1,TCOMBVNCLR,TCOMB_RA1VOR2NF,TCOMB_RA1VOR1NF);
  nand NAND2_6(TCOMBVNODE16,TCOMBVNODE19,TCOMBVNODE16VOR1NF);
  nand NAND2_7(UC_9VZ,UC_9VZVOR1NF,UC_9VUC_0);
  nand NAND2_8(UC_10VZ,UC_10VZVOR1NF,UC_10VUC_0);
  nand NAND2_9(FMLVIINMUXVND1,FMLVIINMUXVOR2NF,FMLVIINMUXVOR1NF);
  nand NAND3_1(TCOMBVNODE3,TCOMBVNODE4,TCOMBVNQB,TCOMBVNQA);
  nand NAND2_10(TESTLVIINMUXVND1,TESTLVIINMUXVOR2NF,TESTLVIINMUXVOR1NF);
  nand NAND2_11(TCOMB_FE,TCOMBVNODE16,TCOMBVNODE14);
  nand NAND2_12(UC_17VUC_0,C2VCO1,UC_17);
  nand NAND2_13(UC_18VUC_0,C2VCO0,UC_18);
  nand NAND2_14(UC_19VUC_0,C2VIINHN,UC_19);
  nand NAND2_15(TCOMB_YA1,TCOMBVNODE16,TCOMBVNODE3);
  nand NAND2_16(UC_17VZ,UC_17VZVOR1NF,UC_17VUC_0);
  nand NAND2_17(UC_18VZ,UC_18VZVOR1NF,UC_18VUC_0);
  nand NAND2_18(UC_19VZ,UC_19VZVOR1NF,UC_19VUC_0);
  nand NAND2_19(C3_Q2VUC_0,C3VCO1,C3_Q2);
  nand NAND2_20(C3_Q1VUC_0,C3VCO0,C3_Q1);
  nand NAND2_21(C3_Q0VUC_0,C3VIINHN,C3_Q0);
  nand NAND2_22(C3_Q2VZ,C3_Q2VZVOR1NF,C3_Q2VUC_0);
  nand NAND2_23(C3_Q1VZ,C3_Q1VZVOR1NF,C3_Q1VUC_0);
  nand NAND2_24(C3_Q0VZ,C3_Q0VZVOR1NF,C3_Q0VUC_0);
  nor NOR3_0(C3VCIIA,C3_Q2,C3_Q1,C3_Q0);
  nor NOR3_1(C1VCIIA,UC_9,UC_10,UC_11);
  nor NOR3_2(C2VCIIA,UC_17,UC_18,UC_19);
  nor NOR2_0(C1_CO,C1VCIIA,UC_12);
  nor NOR3_3(C1VCO2,UC_13,UC_14,UC_15);
  nor NOR2_1(C1VCO1,UC_14,UC_15);
  nor NOR2_2(TCOMBVNODE19,CLRB,TCOMBVNFEL);
  nor NOR4_0(TCOMBVNODE15,CLRB,TCOMBVNFM,TCOMBVNQC,C3_Q1);
  nor NOR2_3(CTST,C1_CO,TESTL);
  nor NOR3_4(UC_11VD,CLRB,UC_11VZ,C1_CO);
  nor NOR4_1(C2VCO2,CTST,C2_QN2,UC_21,UC_22);
  nor NOR3_5(C2VCO1,CTST,UC_21,UC_22);
  nor NOR3_6(C2_CO,C2VCIIA,CTST,UC_20);
  nor NOR2_4(C2VCO0,CTST,UC_22);
  nor NOR4_2(TCOMB_GA2,TCOMB_GA2VAD4NF,TCOMB_GA2VAD3NF,TCOMB_GA2VAD2NF,
    TCOMB_GA2VAD1NF);
  nor NOR2_5(TCOMB_YA2,TCOMBVNODE12,TCOMBVNQA);
  nor NOR2_6(TCOMB_GA1,TCOMBVNODE8,TCOMB_GA1VAD1NF);
  nor NOR3_7(UC_8VD,CLRB,UC_8VZ,C1_CO);
  nor NOR3_8(UC_9VD,CLRB,UC_9VZ,C1_CO);
  nor NOR3_9(UC_10VD,CLRB,UC_10VZ,C1_CO);
  nor NOR4_3(C3VCO2,CO2,UC_24,UC_25,UC_26);
  nor NOR3_10(C3VCO1,CO2,UC_25,UC_26);
  nor NOR3_11(UC_27,C3VCIIA,CO2,UC_23);
  nor NOR2_7(C3VCO0,CO2,UC_26);
  nor NOR3_12(UC_16VD,CLRB,UC_16VZ,C2_CO);
  nor NOR3_13(UC_17VD,CLRB,UC_17VZ,C2_CO);
  nor NOR3_14(UC_18VD,CLRB,UC_18VZ,C2_CO);
  nor NOR3_15(UC_19VD,CLRB,UC_19VZ,C2_CO);
  nor NOR2_8(Y1C,Y1CVAD2NF,Y1CVAD1NF);
  nor NOR2_9(R2C,R2CVAD2NF,R2CVAD1NF);
  nor NOR3_16(C3_Q3VD,CLRB,C3_Q3VZ,UC_27);
  nor NOR3_17(C3_Q2VD,CLRB,C3_Q2VZ,UC_27);
  nor NOR3_18(C3_Q1VD,CLRB,C3_Q1VZ,UC_27);
  nor NOR3_19(C3_Q0VD,CLRB,C3_Q0VZ,UC_27);

endmodule
